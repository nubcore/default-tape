/*
      -- 1 --
     |       |
     6       2
     |       |
      -- 7 --
     |       |
     5       3
     |       |
      -- 4 --
*/

module seg7 (
    input wire [3:0] counter,
    output reg [6:0] segments
);

    always @(*) begin
        case(counter)
            //                7654321
            0:  segments = 7'b1011110; // d
            1:  segments = 7'b1111001; // E
            2:  segments = 7'b1110001; // F
            3:  segments = 7'b1110111; // A
            4:  segments = 7'b0111110; // U
            5:  segments = 7'b0111000; // L
            6:  segments = 7'b1111000; // t
            7:  segments = 7'b0000110; // 1
            8:  segments = 7'b1011011; // 2
            9:  segments = 7'b1001111; // 3
            /*
            0:  segments = 7'b0111111;
            1:  segments = 7'b0000110;
            2:  segments = 7'b1011011;
            3:  segments = 7'b1001111;
            4:  segments = 7'b1100110;
            5:  segments = 7'b1101101;
            6:  segments = 7'b1111101;
            7:  segments = 7'b0000111;
            8:  segments = 7'b1111111;
            9:  segments = 7'b1101111;
            10: segments = 7'b1110111;
            11: segments = 7'b1111100;
            12: segments = 7'b0111001;
            13: segments = 7'b1011110;
            14: segments = 7'b1111001;
            15: segments = 7'b1110001;
            */
	    default:
                segments = 7'b0111111;
        endcase
    end

endmodule
